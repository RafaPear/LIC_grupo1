library ieee;
use ieee.std_logic_1164.all;

entity SerialReceiver is
    port(
        SS
    );
end SerialReceiver;