library ieee;
use ieee.std_logic_1164.all;

entity SLCDC is
    port(
        CLK: in std_logic;
        RESET: in std_logic;
		LCDsel: in std_logic;
        SCLK: in std_logic;
        SDX: in std_logic;
        E: out std_logic;
        D: out std_logic_vector (4 downto 0)
    );
end SLCDC;

architecture arc_slcdc of SLCDC is

component SerialReceiver is
    port(
        SDX: in std_logic;
        SCLK: in std_logic;
        clk_control: in std_logic;
        SS: in std_logic;
        accept: in std_logic;
        RESET: in std_logic;
        D: out std_logic_vector(4 downto 0);
        DX_val: out std_logic
    );
end component;

component LCDDispacher is
    generic(clk_div: natural := 500000);
    port(
        Dval: in std_logic;
        Din: in std_logic_vector(4 downto 0);
        clk: in std_logic;
        Wrl: out std_logic;
        Dout: out std_logic_vector(4 downto 0);
        done: out std_logic
    );
end component;

signal DX_val_temp: std_logic;
signal D_temp: std_logic_vector(4 downto 0);
signal done_temp: std_logic;

begin
USerialReceiver: SerialReceiver
    port map(
        SDX => SDX,
        SCLK => SCLK,
        clk_control => CLK,
        SS => LCDsel,
        accept => done_temp,
        RESET => RESET,
        D => D_temp,
        DX_val => DX_val_temp
    );

UDispacher: LCDDispacher
    port map(
        Dval => DX_val_temp,
        Din => D_temp,
        clk => CLK,
        Wrl => E,
        Dout => D,
        done => done_temp
    );
end arc_slcdc;